----------------------------------------------------------------------------------
-- Company: 
-- Engineer: 
-- 
-- Create Date: 02/15/2025 09:12:12 PM
-- Design Name: 
-- Module Name: Adder_Half - arch_Adder_Half
-- Project Name: 
-- Target Devices: 
-- Tool Versions: 
-- Description: 
-- 
-- Dependencies: 
-- 
-- Revision:
-- Revision 0.01 - File Created
-- Additional Comments:
-- 
----------------------------------------------------------------------------------


library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

-- Uncomment the following library declaration if using
-- arithmetic functions with Signed or Unsigned values
--use IEEE.NUMERIC_STD.ALL;

-- Uncomment the following library declaration if instantiating
-- any Xilinx leaf cells in this code.
--library UNISIM;
--use UNISIM.VComponents.all;

entity Adder_Half is
    Port (
        A : in std_logic;
        B : in std_logic;
        S : out std_logic;
        Cout : out std_logic
    );
end Adder_Half;

architecture arch_Adder_Half of Adder_Half is
    
begin

    S       <= A xor B;
    Cout    <= A and B;

end arch_Adder_Half;